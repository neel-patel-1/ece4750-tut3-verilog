`ifndef ECE4750_TUT3_VERILOG_REGINCR_REG_INCR_V
`define ECE4750_TUT3_VERILOG_REGINCR_REG_INCR_V

module ece4750_tut3_verilog_regincr_Reg_Incr
(
  input logic clk,
  input logic reset,
  input logic [7:0] in_,
  output logic [7:0] out
);

endmodule

`endif // ECE4750_TUT3_VERILOG_REGINCR_REG_INCR_V